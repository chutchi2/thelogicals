** Profile: "SCHEMATIC1-frequ test"  [ C:\Users\Tiffany\Documents\Engineering\ECE4899 - Senior Design\Pspice dummy files\rc test-PSpiceFiles\SCHEMATIC1\frequ test.sim ] 

** Creating circuit file "frequ test.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Tiffany\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC LIN 1000 800Meg 6G
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
