** Profile: "SCHEMATIC1-mc freq"  [ C:\Users\Tiffany\Documents\Engineering\ECE4899 - Senior Design\Pspice dummy files\pfewsma-pspicefiles\schematic1\mc freq.sim ] 

** Creating circuit file "mc freq.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Tiffany\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 100 100 16G
.MC 100 AC V([0]) YMAX LIST OUTPUT ALL SEED=1 
.OPTIONS DISTRIBUTION GAUSS
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
