** Profile: "SCHEMATIC1-mc test"  [ C:\Users\Tiffany\Documents\Engineering\ECE4899 - Senior Design\Pspice dummy files\rc test-PSpiceFiles\SCHEMATIC1\mc test.sim ] 

** Creating circuit file "mc test.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Tiffany\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 2ns 0 
.MC 10 TRAN V([N02150]) YMAX LIST OUTPUT ALL SEED=17366 
.OPTIONS DISTRIBUTION GAUSS
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
